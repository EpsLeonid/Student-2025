package package_settings_V1;
//-----------------------------------------------------------------------------
// Parameter Declaration(s)
//-----------------------------------------------------------------------------
	parameter SIZE_IN_DATA									= 14;
	parameter SIZE_OUT_DATA									= 16;
	parameter SIZE_CNT										= 4;
	parameter DEPTH											= 14;
	parameter k												= 5;
	parameter l												= 8;
	parameter M												= 16;
//-----------------------------------------------------------------------------
endpackage